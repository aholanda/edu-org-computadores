 module hello_world ;
   
   initial begin
      $display ("Alo Mundo");
      #10  $finish;
   end

endmodule 
